Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

Entity Cont4_mod10 is
    PORT(RST  : in std_logic;
         CLK  : in std_logic;
         EN   : in std_logic;
         CLR  : in std_logic;
         Q    : out unsigned(3 downto 0);
         COUT : out std_logic
    );
end entity;

Architecture X of Cont4_mod10 is
    Signal CONT: unsigned (3 downto 0) := (others => '0');
    Begin
    Process (CLK, RST)
    Begin
        If RST = '1' then
            CONT <= "0000";
        Elsif CLK' event and CLK = '1' then
            If CLR = '1'then
                CONT <= "0000";
            Else
                If EN = '1' then
                    If CONT = "1001" then
                        CONT <= (others => '0');
                    Else
                        CONT <= CONT + 1;
                    End IF;
                End If;
            End If;
        End If;
    End process;
    Q <= CONT;
    COUT <= '1' when (EN='1' and CONT = "1001") else '0';
End architecture;
